----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:52:08 11/16/2023 
-- Design Name: 
-- Module Name:    new_sbox3 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
	Library UNISIM;
	use UNISIM.vcomponents.all;
		use std.textio.all;
	use ieee.std_logic_textio.all;

entity new_sbox3 is
port(
      DO : out  std_logic_vector(31 downto 0);      -- 32-bit Data Output
      DOP : out  std_logic_vector(3 downto 0);    -- 4-bit parity Output
      ADDR : in integer;   -- 9-bit Address Input
      CLK : in std_logic;   -- Clock
      DI : in std_logic_vector(31 downto 0);      -- 32-bit Data Input
      DIP :in std_logic_vector(3 downto 0);  -- 4-bit parity Input
      EN : in std_logic;     -- RAM Enable Input
      SSR :in std_logic;   -- Synchronous Set/Reset Input
      WE : in std_logic
);
end new_sbox3;

architecture Behavioral of new_sbox3 is
signal address : std_logic_vector(8 downto 0);

begin


address <= std_logic_vector(to_unsigned(addr,9));
------------------------sbox 3----------------------------------------------------------

RAMB16_S36_inst : RAMB16_S36
   generic map (
      INIT => X"000000000",  --  Value of output RAM registers at startup
      SRVAL => X"000000000", --  Output value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Address 0 to 127
      INIT_00 => X"d4a20068bcf46b2e7602d4f7411520f794692934f64c261c948140f7e93d5a68",
      INIT_01 => X"bf8b884014214f74972445461e39f62e500061af43b7d4b73320f46ad4082471",
      INIT_02 => X"31cb85047fac6dd003bd9785bfbc09ec66a02f4570f4ddd396b591af4d95fc1d",
      INIT_03 => X"e9b66dfb0a2c86da530429f428507825abca0a9ada2547e655fd394196eb27b3",
      INIT_04 => X"7af4d6b6b58ce006e887ad8c4f3ffea227a18dee680ec0a4d748690068dc1462",
      INIT_05 => X"3b124e8bee39d7abd9f385b920fe9e35406b2a42ce78a399d3375fecaace1e7c",
      INIT_06 => X"ca7820fb6841e7f7dd5b43323a6efa74eae397b226a366314b6d18561dc9faf7",
      INIT_07 => X"d096954bfe6ba9b720838d8755533a3aba489527454056acd8feb397fb0af54e",
      INIT_08 => X"9029317c5ef47e1c3f3125f9a62a4a5699e1db33cca92963a1159a5855a867bc",
      INIT_09 => X"c70f86dc48c1133fe4c66d2295c1154805282ce380bb155c04272f70fdf8e802",
      INIT_0A => X"41113564f2bcc18fd59bc0d1325f51eb5d886e17404779a441041f0f07f9c9ee",
      INIT_0B => X"cad18115af664fd102e1329e0e12b4c21f636c1bdff8e8a3602a9c60257b7834",
      INIT_0C => X"2da2f728de720c8ce6ba0d9985b2a20eeebeb9223b240b62333e92e16b2395e0",
      INIT_0D => X"f33e8d1ec39dfd27877d48fa5449a36fe7ccf5f0647d086295b794fdd0127845",
      INIT_0E => X"db6e6b0d991be14ca1ebddf8a812dc60f4f8fd373a6f6eab992eff740a476341",
      INIT_0F => X"690fed0bb5390f92cc00ffa3f1290dc7dcd0e8042765d43b6d672c37c67b5510",
      -- Address 128 to 255
      INIT_10 => X"763bd6eb7b9479bf515bad24bb132f88d9155ea3a091cf0bcedb7d9c667b9ffb",
      INIT_11 => X"782ef11c12754cccc66a2b3b6842ada7f42e312d8026e297cc11597937392eb3",
      INIT_12 => X"e2e1c3c93d25bdd811caedfa1a6b10184bfb635006a1bbe6b79251e76a124237",
      INIT_13 => X"64e4c3febebfe988da86a85f64af674ed5abea2ad90cec6e0a12138644421659",
      INIT_14 => X"d736fccc7745ae04f6381fb0d1fd83466003604d60787bf8f0f7c0869dbc8057",
      INIT_15 => X"bf582e6155464299bde8ae2477a057be3c005e5fb0804187f01eab7183426b33",
      INIT_16 => X"46fcd9b9b475f255c8b38e745366f9c38789bdc2f474ef38f2ddfda24e58f48f",
      INIT_17 => X"c902de4c8cd5559120b45770466e598e915f95e2846a0e798b1ddf847aeb2661",
      INIT_18 => X"c4324633662d09a1e0a9dc09b77f19b67574a99e11a86248bb8205d0b90bace1",
      INIT_19 => X"2868f169a186f20f0ba5a4df1ab93d1d1d6efe104a99a02509f0be8ce85a1f02",
      INIT_1A => X"0de6d027a002b5c4a70683fa50115e014fcd7f52a1e2ce9b573906fedcb7da83",
      INIT_1B => X"30dc7d62006058aac0f586e0f0177a2861a806b5c3604c06773f86419af88c27",
      INIT_1C => X"ce591d76ebfc7da190bcb6debbcbee56c2c2163453c2dd942338ea6311e69ed7",
      INIT_1D => X"d39eb8fc1ac15bb4724d9db986e3725f7c927c2439720a3d4b7c01886f05e409",
      INIT_1E => X"6c51133ca28514d9b161e6f81e50ef5e4dad0fc4d83d7cd308fca5b5ed545578",
      INIT_1F => X"406000e0670efa8e92638212d79a3234ddc6c837362abfce56e14ec46fd5c7e7",
      -- Address 256 to 383
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 384 to 511
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Address 0 to 127
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 128 to 255
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 256 to 383
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 384 to 511
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO => DO,      -- 32-bit Data Output
      DOP => DOP,    -- 4-bit parity Output
      ADDR => address,  -- 9-bit Address Input
      CLK => CLK,    -- Clock
      DI => DI,      -- 32-bit Data Input
      DIP => DIP,    -- 4-bit parity Input
      EN => EN,      -- RAM Enable Input
      SSR => SSR,    -- Synchronous Set/Reset Input
      WE => WE       -- Write Enable Input
   );



end Behavioral;

