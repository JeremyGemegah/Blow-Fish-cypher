----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:52:26 11/16/2023 
-- Design Name: 
-- Module Name:    new_sbox4 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
	Library UNISIM;
	use UNISIM.vcomponents.all;
		use std.textio.all;
	use ieee.std_logic_textio.all;


entity new_sbox4 is
port(
      DO : out  std_logic_vector(31 downto 0);      -- 32-bit Data Output
      DOP : out  std_logic_vector(3 downto 0);    -- 4-bit parity Output
      ADDR : in  integer;   -- 9-bit Address Input
      CLK : in std_logic;   -- Clock
      DI : in std_logic_vector(31 downto 0);      -- 32-bit Data Input
      DIP :in std_logic_vector(3 downto 0);  -- 4-bit parity Input
      EN : in std_logic;     -- RAM Enable Input
      SSR :in std_logic;   -- Synchronous Set/Reset Input
      WE : in std_logic
);
end new_sbox4;

architecture Behavioral of new_sbox4 is
signal address: std_logic_vector(8 downto 0);

begin

address <= std_logic_vector(to_unsigned(addr,9));

---------------------------------sbox 4 -------------------------------------------------------

RAMB16_S36_inst : RAMB16_S36
   generic map (
      INIT => X"000000000",  --  Value of output RAM registers at startup
      SRVAL => X"000000000", --  Output value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Address 0 to 127
      INIT_00 => X"99bc9bbed38227404fa337425cb0679e5ac52d1babc27737d3faf5cf3a39ce37",
      INIT_01 => X"6a366eb4b26eb1be21a19045b78c1b6bc700c47bd62d1c7ebf0f7315d5118e9d",
      INIT_02 => X"4cd04dc6d5730a1d468dde7d530ff8ee6549c2c8c6a376d2bc946e795748ab2f",
      INIT_03 => X"9a86ee2263ef8ce26a2d519aa1fad5f0be5ee304ac9526e8a9ba46502939bbdb",
      INIT_04 => X"ba645bd68fe515509be96a4d83c061ba9cf2d0a4a51e03aa43242ef6c089c2b8",
      INIT_05 => X"77fa0a593f046f69f752f7dac72fefd3ef5562e94ba99586a73a3ae12826a2f9",
      INIT_06 => X"022b8b512cf0b7d99e34d797e990fd5a3b3ee5939b09e6ad87b0860180e4a915",
      INIT_07 => X"5a88f54c5ad6b472adf2b89b1f9f25cf7c7d2d28d1cf3ed6017da67d96d5ac3a",
      INIT_08 => X"79132e28f8d56629283b57cce8d3c48ded93fa9b47b0acfde019a5e6e029ac71",
      INIT_09 => X"0564f0bd03a1612588f46dba15056dd4e3d35e8cf7960e44ed756055785f0191",
      INIT_0A => X"26dcf319f59c66fb1e6321f51b3f6d9ba93a072a97271aec3c9057a2c3eb9e15",
      INIT_0B => X"ccad925fabcc5167c20ad9f8285177118aba3cbb03563482b155fdf57533d928",
      INIT_0C => X"774fbe325121ce64fb3e7bceea7a90c29320f991379d58623830dc8e4de81751",
      INIT_0D => X"0907216669852dfddd6db224a2ae08106413e68048de5369c3293d46a8b6e37e",
      INIT_0E => X"6bb4e3bbccd2017f1b588d405bbef7dd1c20c8ae586cdecf6445c0ddb39a460a",
      INIT_0F => X"bf3c6f478d6612aefa6484bb72eacea8bcb4cdd53e350a443a59ff45dda26a7e",
      -- Address 128 to 255
      INIT_10 => X"af537d5df8721671e75b1357740e0d8df64e6370aec2771b542f5d9ed29be463",
      INIT_11 => X"ce6ea04806b89fb495983a1de1b004280115af8434d2466a4eb4e2cc4040cb08",
      INIT_12 => X"344525bdbb3a792be7933fdc611560b1277227f8011a1d4b3520ab826f3f3b82",
      INIT_13 => X"a1e8aac7cf0111c3bcc7d1f6e01cc87ea01fbac92f32c9b751ce794ba08839e1",
      INIT_14 => X"e0b12b4f8df9317cc69136670339c32ad50ada38d0dadecbd44fbd9a1a908749",
      INIT_15 => X"9b9415250f91fc7115e6fc2abf97222c27d9459cf2d519ff43f5bb3af79e59b7",
      INIT_16 => X"cb03a44210d25065e3056a0cb6c1075e12baa8d1c2a86459ceb69cebfae59361",
      INIT_17 => X"8971f21ed3a0342be0d392df9f1f95323278e9644c98a0be1698db3be0ec6e0e",
      INIT_18 => X"0fe3f11de60b6f479b992f2edf359f8dc37632d8c5be71204ba3348c1b0a7441",
      INIT_19 => X"f6fb2299848fd2c5fd2c1d051618b166cd3e7e6fce6279cf1edad891e54cda54",
      INIT_1A => X"88d273cc6e1636975a75ebb5acf0816256cccd0293a83531a6327623f523f357",
      INIT_1B => X"c3f27b9a45e1d006327a140ae6c6c7bd71c656144c50901b81b949d0de966292",
      INIT_1C => X"cd769c2bb6cbcf7cb20402227112690535bdd2f6bb25bfe262a80f00c9aa53fd",
      INIT_1D => X"2075606077afa1c5f746ce76ba38209c2547adf038abbd601640e3d353113ec0",
      INIT_1E => X"d6ebe1f901c36ae402fb8a8c1948c25c4cf9aa7e7aaaf9b08ae88dd885cbfe4e",
      INIT_1F => X"3ac372e6578fdfe3ce77e25bb74e6132c208e69f3f09252da65cdea090d4f869",
      -- Address 256 to 383
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 384 to 511
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Address 0 to 127
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 128 to 255
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 256 to 383
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 384 to 511
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO => DO,      -- 32-bit Data Output
      DOP => DOP,    -- 4-bit parity Output
      ADDR => address,  -- 9-bit Address Input
      CLK => CLK,    -- Clock
      DI => DI,      -- 32-bit Data Input
      DIP => DIP,    -- 4-bit parity Input
      EN => EN,      -- RAM Enable Input
      SSR => SSR,    -- Synchronous Set/Reset Input
      WE => WE       -- Write Enable Input
   );

end Behavioral;

